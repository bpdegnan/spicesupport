* Transmission gate characterization
* Standard t-gate vs m=2 vs mulid0=2

* Include the PDK models
.lib $SPICE_LIB/sky130.lib.spice tt

* Include abstract device definitions
.include devices.cir

* Supply
Vdd vdd 0 DC 1.8

* Shared sweep voltage
Vcm cm 0 DC 0

* Standard transmission gate (m=1)
Xn1 in1 vdd cm 0 abnmos
Xp1 in1 0 cm vdd abpmos
Vds1 in1 cm DC 0.025

* Transmission gate with m=2
Xn2 in2 vdd cm 0 abnmos m=2
Xp2 in2 0 cm vdd abpmos m=2
Vds2 in2 cm DC 0.025

* Transmission gate with mulid0=2
Xn3 in3 vdd cm 0 abnmos mulid0=2
Xp3 in3 0 cm vdd abpmos mulid0=2
Vds3 in3 cm DC 0.025

.control
    dc Vcm 0 1.8 0.001
    set wr_vecnames
    set wr_singlescale
    wrdata tgatedc.csv v(cm) i(Vds1) i(Vds2) i(Vds3)
    echo "Done"
.endc

.end