* NFET Transient gate sweep - HSPICE version
* Gate ramps from 0V to VDD over 1ms
* Measures all terminal currents: gate, drain, source, bulk
* For comparing behavior across different systems/configurations

* HSPICE options
* post=2 should give ASCII
* .option post=2
* RUNLVL=6 as explicit options
.option method=gear
* bypass of 2 is for MOSFETS, 0 calculate everything
.option bypass=0
.option accurate=1
.option reltol=1e-5
.option abstol=1e-15
.option vntol=1e-7
.option absi=1e-15
.option absmos=1e-15
.option lvltim=3 
.option dvdt=2
* trtol is a bit of a mystery as it's used as an error estimator.  1 is unity
.option trtol=1  

* pivot/matrix issues for pivot too large warning
.option gmin=1e-15
.option gmindc=1e-15
.option pivot=13
.option pivrel=1e-3


*more transient options to try to fix wave
.option delmax=1e-6
.option bytol=1e-6

* Include the HSPICE-compatible PDK library
.lib '../sky130.l' tt
.include '../devices_hspice.cir'

* Parameters
.param VDD_VAL=1.8

* Supply
Vdd vdd 0 DC VDD_VAL

* Gate voltage ramp with current sensing (0 to 1.8V over 1ms)
Vg ng_int 0 PWL(0 0 1m VDD_VAL)
Vg_sense ng_int ng DC 0

* Drain at VDD with current sensing
Vd vdd nd_int DC 0
Vd_sense nd_int nd DC 0

* Source at ground with current sensing
Vs_sense ns 0 DC 0

* Bulk at ground with current sensing
Vb_sense nb 0 DC 0

* NFET: drain, gate, source, bulk
Xnmos nd ng ns nb abnmos

* Transient analysis: 1ms with some timestep.  
.tran 1u 1m

* Output currents
.print tran v(ng) i(Vg_sense) i(Vd_sense) i(Vs_sense) i(Vb_sense)

.end
