* PFET gate sweep at two drain voltages - HSPICE version

* HSPICE options
.option post accurate

* Include the HSPICE-compatible PDK library
.lib '../../sky130.l' tt
.include '../../devices_hspice.cir'

* Supply
Vdd vdd 0 DC 1.8

* PFET at Vd=0V (saturation, |Vds|=1.8V)
Xpmos_sat pd_sat ng vdd vdd abpmos
Vp_sat pd_sat 0 DC 0

* PFET at Vd=1.7V (linear, |Vds|=100mV)
Xpmos_lin pd_lin ng vdd vdd abpmos
Vp_lin pd_lin 0 DC 1.7

* Shared gate
Vg ng 0 DC 0

* DC sweep of gate voltage
.dc Vg 0 1.8 0.001

* Output currents
.print dc v(ng) i(Vp_sat) i(Vp_lin)

.end
