* PFET gate sweep at two drain voltages - ngspice version

* Include the PDK models
.lib $SPICE_LIB/sky130.lib.spice tt

* Include abstract device definitions
.include ../../devices_ngspice.cir

* Supply
Vdd vdd 0 DC 1.8

* PFET at Vd=0V (saturation, |Vds|=1.8V)
Xpmos_sat pd_sat ng vdd vdd abpmos
Vp_sat pd_sat 0 DC 0

* PFET at Vd=1.7V (linear, |Vds|=100mV)
Xpmos_lin pd_lin ng vdd vdd abpmos
Vp_lin pd_lin 0 DC 1.7

* Shared gate
Vg ng 0 DC 0

.control
    dc Vg 0 1.8 0.001
    set wr_vecnames
    set wr_singlescale
    wrdata pfet_ngspice.csv v(ng) i(Vp_sat) i(Vp_lin)
    echo "Done"
.endc

.end
