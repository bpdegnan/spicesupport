* Common source amplifier - NMOS and PMOS versions


* Include the PDK models
.lib $SPICE_LIB/sky130.lib.spice tt

* Include abstract device definitions
.include devices.cir

* Supply
Vdd vdd 0 DC 1.8

* NMOS: Bottom nFET as bias, top nFET as input
* 100mV bias
Xn_bias1 voutn1 nbias1 0 0 abnmos
Vbias_n1 nbias1 0 DC 0.1
Xn_in1 vdd in voutn1 0 abnmos

* 200mV bias
Xn_bias2 voutn2 nbias2 0 0 abnmos
Vbias_n2 nbias2 0 DC 0.2
Xn_in2 vdd in voutn2 0 abnmos

* PMOS: Top pFET as bias, bottom pFET as input
* 100mV bias (1.7V = VDD - 100mV)
Xp_bias1 voutp1 pbias1 vdd vdd abpmos
Vbias_p1 pbias1 0 DC 1.7
Xp_in1 0 in voutp1 vdd abpmos

* 200mV bias (1.6V = VDD - 200mV)
Xp_bias2 voutp2 pbias2 vdd vdd abpmos
Vbias_p2 pbias2 0 DC 1.6
Xp_in2 0 in voutp2 vdd abpmos

* Input sweep
Vin in 0 DC 0

.control
    dc Vin 0 1.8 0.001
    set wr_vecnames
    set wr_singlescale
    wrdata commonsource.csv v(in) v(voutn1) v(voutn2) v(voutp1) v(voutp2)
    echo "Done"
.endc

.end