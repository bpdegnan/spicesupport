* Abstract devices for HSPICE with SkyWater 130nm PDK
* These bypass the ngspice-specific subcircuits

* NMOS transistor subcircuit definition
.subckt abnmos D G S B l=0.15u w=1u
M1 D G S B sky130_fd_pr__nfet_01v8 l=l w=w
.ends abnmos

* PMOS transistor subcircuit definition
.subckt abpmos D G S B l=0.15u w=1u
M1 D G S B sky130_fd_pr__pfet_01v8 l=l w=w
.ends abpmos